library verilog;
use verilog.vl_types.all;
entity fvc_tst is
end fvc_tst;
