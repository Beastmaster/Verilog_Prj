-- megafunction wizard: %Serial Flash Loader%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altserial_flash_loader 

-- ============================================================
-- File Name: ok.vhd
-- Megafunction Name(s):
-- 			altserial_flash_loader
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.0 Build 235 06/17/2009 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY ok IS
	PORT
	(
		asdo_in		: IN STD_LOGIC ;
		asmi_access_granted		: IN STD_LOGIC ;
		dclk_in		: IN STD_LOGIC ;
		ncso_in		: IN STD_LOGIC ;
		noe_in		: IN STD_LOGIC ;
		asmi_access_request		: OUT STD_LOGIC ;
		data0_out		: OUT STD_LOGIC 
	);
END ok;


ARCHITECTURE SYN OF ok IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT altserial_flash_loader
	GENERIC (
		enable_shared_access		: STRING;
		enhanced_mode		: NATURAL;
		intended_device_family		: STRING;
		lpm_type		: STRING
	);
	PORT (
			scein	: IN STD_LOGIC ;
			dclkin	: IN STD_LOGIC ;
			data0out	: OUT STD_LOGIC ;
			sdoin	: IN STD_LOGIC ;
			asmi_access_granted	: IN STD_LOGIC ;
			asmi_access_request	: OUT STD_LOGIC ;
			noe	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	data0_out    <= sub_wire0;
	asmi_access_request    <= sub_wire1;

	altserial_flash_loader_component : altserial_flash_loader
	GENERIC MAP (
		enable_shared_access => "ON",
		enhanced_mode => 1,
		intended_device_family => "Cyclone II",
		lpm_type => "altserial_flash_loader"
	)
	PORT MAP (
		scein => ncso_in,
		dclkin => dclk_in,
		sdoin => asdo_in,
		asmi_access_granted => asmi_access_granted,
		noe => noe_in,
		data0out => sub_wire0,
		asmi_access_request => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ENABLE_SHARED_ACCESS STRING "ON"
-- Retrieval info: CONSTANT: ENHANCED_MODE NUMERIC "1"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: USED_PORT: asdo_in 0 0 0 0 INPUT NODEFVAL "asdo_in"
-- Retrieval info: USED_PORT: asmi_access_granted 0 0 0 0 INPUT NODEFVAL "asmi_access_granted"
-- Retrieval info: USED_PORT: asmi_access_request 0 0 0 0 OUTPUT NODEFVAL "asmi_access_request"
-- Retrieval info: USED_PORT: data0_out 0 0 0 0 OUTPUT NODEFVAL "data0_out"
-- Retrieval info: USED_PORT: dclk_in 0 0 0 0 INPUT NODEFVAL "dclk_in"
-- Retrieval info: USED_PORT: ncso_in 0 0 0 0 INPUT NODEFVAL "ncso_in"
-- Retrieval info: USED_PORT: noe_in 0 0 0 0 INPUT NODEFVAL "noe_in"
-- Retrieval info: CONNECT: @sdoin 0 0 0 0 asdo_in 0 0 0 0
-- Retrieval info: CONNECT: asmi_access_request 0 0 0 0 @asmi_access_request 0 0 0 0
-- Retrieval info: CONNECT: @dclkin 0 0 0 0 dclk_in 0 0 0 0
-- Retrieval info: CONNECT: @scein 0 0 0 0 ncso_in 0 0 0 0
-- Retrieval info: CONNECT: @noe 0 0 0 0 noe_in 0 0 0 0
-- Retrieval info: CONNECT: @asmi_access_granted 0 0 0 0 asmi_access_granted 0 0 0 0
-- Retrieval info: CONNECT: data0_out 0 0 0 0 @data0out 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ok.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ok.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ok.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ok.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ok_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
