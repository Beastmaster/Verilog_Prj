module stopwatch(EN,CP,cntH,cntL);



endmodule 